package uart_pkg;

	`include "uart_transaction.sv"
	`include "uart_generator.sv"
	`include "uart_driver.sv"
	`include "uart_monitor.sv"
	`include "uart_scoreboard.sv"
	`include "uart_environment.sv"
	
endpackage